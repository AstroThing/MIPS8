`timescale 1ns / 1ps

module CPU(
    input clk,
	 output reg [7:0] data
    );


endmodule
