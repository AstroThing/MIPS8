`timescale 1ns / 1ps

module Main(
    input clk
    );

	CPU cpu(clk);
endmodule
