`timescale 1ns / 1ps

module CPU(
    input clk
    );

reg [7:0] PC;

endmodule
